
        
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;
-- use IEEE.fixed_pkg.all;

        package dtypes is
            type int_array is array (0 to 600) of integer;
        end package;

        
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;
-- use IEEE.fixed_pkg.all;

        
library work;       -- Default package name
use work.config.all;

        use work.dtypes.all;
        
        entity sigmoid is
            port (
                clk    : in std_logic;
                en     : in std_logic;
                num    : in integer;
                result : out integer;
                done   : out std_logic
            );
        end sigmoid;
        

        architecture Behavioral of sigmoid is
        begin

            process(clk)
            variable sigm : int_array := (268,270,272,274,276,278,280,282,284,286,289,291,293,295,297,299,301,303,305,307,310,312,314,316,318,320,323,325,327,329,331,334,336,338,340,342,345,347,349,352,354,356,358,361,363,365,368,370,372,375,377,379,382,384,386,389,391,394,396,398,401,403,406,408,410,413,415,418,420,423,425,428,430,432,435,437,440,442,445,447,450,452,455,457,460,462,465,467,470,472,475,477,480,482,485,487,490,492,495,497,500,502,504,507,509,512,514,517,519,522,524,527,529,532,534,537,539,542,544,547,549,552,554,557,559,562,564,567,569,571,574,576,579,581,584,586,589,591,593,596,598,601,603,605,608,610,613,615,617,620,622,624,627,629,631,634,636,638,641,643,645,647,650,652,654,657,659,661,663,665,668,670,672,674,676,679,681,683,685,687,689,692,694,696,698,700,702,704,706,708,710,713,715,717,719,721,723,725,727,729,731,733,734,736,738,740,742,744,746,748,750,752,753,755,757,759,761,763,764,766,768,770,772,773,775,777,779,780,782,784,785,787,789,790,792,794,795,797,798,800,802,803,805,806,808,809,811,813,814,816,817,819,820,822,823,824,826,827,829,830,832,833,834,836,837,838,840,841,842,844,845,846,848,849,850,851,853,854,855,856,858,859,860,861,862,864,865,866,867,868,869,871,872,873,874,875,876,877,878,879,880,881,882,883,884,885,886,887,888,889,890,891,892,893,894,895,896,897,898,899,900,901,902,902,903,904,905,906,907,908,908,909,910,911,912,912,913,914,915,916,916,917,918,919,919,920,921,922,922,923,924,924,925,926,926,927,928,928,929,930,930,931,932,932,933,934,934,935,935,936,937,937,938,938,939,939,940,941,941,942,942,943,943,944,944,945,945,946,946,947,947,948,948,949,949,950,950,951,951,952,952,953,953,953,954,954,955,955,956,956,956,957,957,958,958,958,959,959,960,960,960,961,961,961,962,962,963,963,963,964,964,964,965,965,965,966,966,966,967,967,967,968,968,968,968,969,969,969,970,970,970,970,971,971,971,972,972,972,972,973,973,973,973,974,974,974,974,975,975,975,975,976,976,976,976,977,977,977,977,977,978,978,978,978,978,979,979,979,979,979,980,980,980,980,980,981,981,981,981,981,982,982,982,982,982,982,983,983,983,983,983,983,984,984,984,984,984,984,984,985,985,985,985,985,985,985,986,986,986,986,986,986,986,987,987,987,987,987,987,987,987,987,988,988,988,988,988,988,988,988,989,989,989,989,989,989,989,989,989,989,990,990,990,990,990,990,990,990,990,990,990,991,991,991,991,991,991,991,991,991,991,991,991,992,992,992,992,992,992,992,992,992,992,992,992,992,993,993,993,993,993);
            begin

                if rising_edge(clk) then
                    if EN = '1' and num > -100.0 and num < 6000 then
                        result <= sigm((100) + num/10); -- take note of precision if 0.1 leave as is if 0.01 divide by 1
                        done <= '1';
                    else
                        done <= '0';
                    end if;
                end if;
            end process;
        end behavioral;
        