
        
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;
-- use IEEE.fixed_pkg.all;

        package dtypes is
            type int_array is array (0 to 600) of integer;
        end package;

        
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;
-- use IEEE.fixed_pkg.all;

        
library work;       -- Default package name
use work.config.all;

        use work.dtypes.all;
        
        entity tanh_activation is
            port (
                clk    : in std_logic;
                en     : in std_logic;
                num    : in integer;
                result : out integer;
                done   : out std_logic
            );
        end tanh_activation;
        

        architecture Behavioral of tanh_activation is
        begin

            process(clk)
            variable tanh : int_array := (-761,-757,-753,-748,-744,-739,-735,-730,-725,-721,-716,-711,-706,-701,-696,-691,-685,-680,-675,-669,-664,-658,-652,-646,-641,-635,-629,-623,-616,-610,-604,-597,-591,-584,-578,-571,-564,-558,-551,-544,-537,-529,-522,-515,-507,-500,-492,-485,-477,-469,-462,-454,-446,-438,-430,-421,-413,-405,-396,-388,-379,-371,-362,-353,-345,-336,-327,-318,-309,-300,-291,-282,-272,-263,-254,-244,-235,-226,-216,-206,-197,-187,-178,-168,-158,-148,-139,-129,-119,-109,-99,-89,-79,-69,-59,-49,-39,-29,-19,-9,0,9,19,29,39,49,59,69,79,89,99,109,119,129,139,148,158,168,178,187,197,206,216,226,235,244,254,263,272,282,291,300,309,318,327,336,345,353,362,371,379,388,396,405,413,421,430,438,446,454,462,469,477,485,492,500,507,515,522,529,537,544,551,558,564,571,578,584,591,597,604,610,616,623,629,635,641,646,652,658,664,669,675,680,685,691,696,701,706,711,716,721,725,730,735,739,744,748,753,757,761,765,769,773,777,781,785,789,793,796,800,804,807,811,814,817,821,824,827,830,833,836,839,842,845,848,851,853,856,859,861,864,866,869,871,874,876,878,880,883,885,887,889,891,893,895,897,899,901,903,905,906,908,910,912,913,915,917,918,920,921,923,924,926,927,928,930,931,932,934,935,936,937,939,940,941,942,943,944,945,946,947,948,949,950,951,952,953,954,955,956,957,957,958,959,960,961,961,962,963,964,964,965,966,966,967,968,968,969,969,970,971,971,972,972,973,973,974,974,975,975,976,976,977,977,978,978,978,979,979,980,980,980,981,981,981,982,982,983,983,983,983,984,984,984,985,985,985,986,986,986,986,987,987,987,987,988,988,988,988,989,989,989,989,989,990,990,990,990,990,991,991,991,991,991,991,992,992,992,992,992,992,992,993,993,993,993,993,993,993,993,994,994,994,994,994,994,994,994,994,995,995,995,995,995,995,995,995,995,995,995,996,996,996,996,996,996,996,996,996,996,996,996,996,996,996,997,997,997,997,997,997,997,997,997,997,997,997,997,997,997,997,997,997,997,997,998,998,998,998,998,998,998,998,998,998,998,998,998,998,998,998,998,998,998,998,998,998,998,998,998,998,998,998,998,998,998,998,998,998,998,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999,999);
            begin

                if rising_edge(clk) then
                    if EN = '1' then
                        if num > -1000 and num < 6000 then
                            result <= sigm((100) + num/10); -- take note of precision if 0.1 leave as is if 0.01 divide by 1
                            done <= '1';
                        else
                            result <= 0;
                            done <= '1';
                        end if;
                    else
                        done <= '0';
                    end if;
                end if;
            end process;
        end behavioral;
        